library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.wishbone_pkg.all;


entity blinky is

    port(
    
    -- these two sys signal come from SysCon
    s_clk_sys_i       : in std_ulogic;
    s_rst_sys_n_i       : in std_ulogic;


    t_wb_out          : out t_wishbone_slave_out;
      -- type t_wishbone_slave_out is record
      -- ack   : std_logic;
      -- err   : std_logic;
      -- rty   : std_logic;
      -- stall : std_logic;
      -- dat   : t_wishbone_data;
      -- end record t_wishbone_slave_out;

    t_wb_in            : in  t_wishbone_slave_in;
      --type t_wishbone_slave_in is record
      --cyc : std_logic;
      --stb : std_logic;
      --adr : t_wishbone_address;
      --sel : t_wishbone_byte_select;
      --we  : std_logic;
      --dat : t_wishbone_data;
      --end record t_wishbone_slave_in;

    s_led_o           : out std_logic
    );

end entity;

architecture blinky_arch of blinky is

  --signal s_rst_sys_n        : std_logic := '0';
  signal s_led_state        : std_logic := '0';
  signal s_stall_state      : std_logic := '0';

  --signal s_led_freq_ctl     : std_logic := '0';
  --signal s_count            : integer   :=  1;
  --signal s_compare_to       : integer   :=  1;

  --signal  s_blinky_mode_v   : std_logic_vector(2 downto 0);

  --constant s_blinky_mode_A  : std_logic_vector(2 downto 0) := "000";
  --constant s_blinky_mode_B  : std_logic_vector(2 downto 0) := "001";
  --constant s_blinky_mode_C  : std_logic_vector(2 downto 0) := "100";

begin
  
  --  for now no errors, no stalling
  t_wb_out.err    <= '0';
  t_wb_out.stall  <= s_stall_state;
  t_wb_out.rty    <= '0';

  t_wb_out.ack <= t_wb_in.stb and t_wb_in.cyc;

  s_led_o <= s_led_state;
  --s_led_o <= s_led_state and s_led_freq_ctl;

  -- single read write cycle
  p_wb_read_write: process(s_clk_sys_i, s_rst_sys_n_i)

  begin

  if rising_edge(s_clk_sys_i) then

    -- RESET
    -- reset is active low
    if (s_rst_sys_n_i = '0') then
      if rising_edge(s_clk_sys_i) then
      -- all wishbone interfaces must initialize on the rising clock 
      -- after reset was called

      -- RESET
      t_wb_out.dat    <= (others => '0');

      s_led_state     <= '0';
      s_stall_state   <= '0';

      --s_blinky_mode_v   <= (others => '0');
      --s_led_freq_ctl  <= '1';
      --s_count         <=  1;
      --s_compare_to    <=  15; --15000
      end if; --rising_edge(s_clk_sys_i)

      -- END t_wb_in.stb = '1' and t_wb_in.cyc = '1' and t_wb_in.we = '1'

    -- WRITE
    elsif t_wb_in.stb = '1' and t_wb_in.cyc = '1' and t_wb_in.we = '1' then

      s_led_state        <= t_wb_in.dat(0);
      
      -- END WRITE
      -- END t_wb_in.stb = '1' and t_wb_in.cyc = '1' and t_wb_in.we = '1'
  
    -- READ
    elsif t_wb_in.stb = '1' and t_wb_in.cyc = '1' and t_wb_in.we = '0' then
      
      t_wb_out.dat(0) <= s_led_state;
      
      -- END READ
      -- END t_wb_in.stb = '1' and t_wb_in.cyc = '1' and t_wb_in.we = '0'


    end if;

  -- END rising_edge(s_clk_sys_i)
  end if;

  end process;
            
end blinky_arch;